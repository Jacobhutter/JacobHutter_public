library verilog;
use verilog.vl_types.all;
entity bp_sv_unit is
end bp_sv_unit;
