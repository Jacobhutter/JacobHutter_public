module rotation(input Clk,Reset,rotate_enable,
					 input [9:0] square1x,square1y,square2x,square2y,square3x,square3y,square4x,square4y,
					 input [3:0] shape,
					 output square1);

endmodule
