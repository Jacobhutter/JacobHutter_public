library verilog;
use verilog.vl_types.all;
entity mem_control_sv_unit is
end mem_control_sv_unit;
