library verilog;
use verilog.vl_types.all;
entity tagwrite_sv_unit is
end tagwrite_sv_unit;
