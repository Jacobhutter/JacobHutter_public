library verilog;
use verilog.vl_types.all;
entity wishbone_interface_sv_unit is
end wishbone_interface_sv_unit;
