library verilog;
use verilog.vl_types.all;
entity evictbuffer is
end evictbuffer;
