library verilog;
use verilog.vl_types.all;
entity tagchecker4_sv_unit is
end tagchecker4_sv_unit;
