library verilog;
use verilog.vl_types.all;
entity ebdatapath_sv_unit is
end ebdatapath_sv_unit;
