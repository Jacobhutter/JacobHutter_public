library verilog;
use verilog.vl_types.all;
entity wordswap_sv_unit is
end wordswap_sv_unit;
