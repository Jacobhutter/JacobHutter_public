library verilog;
use verilog.vl_types.all;
entity tagchecker_sv_unit is
end tagchecker_sv_unit;
