library verilog;
use verilog.vl_types.all;
entity mem_controller_sv_unit is
end mem_controller_sv_unit;
