library verilog;
use verilog.vl_types.all;
entity cachelru4_sv_unit is
end cachelru4_sv_unit;
