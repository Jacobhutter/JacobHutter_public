library verilog;
use verilog.vl_types.all;
entity selectway4_sv_unit is
end selectway4_sv_unit;
