library verilog;
use verilog.vl_types.all;
entity interconnect is
end interconnect;
