library verilog;
use verilog.vl_types.all;
entity swapaddress_sv_unit is
end swapaddress_sv_unit;
