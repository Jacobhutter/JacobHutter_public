import lc3b_types::*;

module cache
(
    input clk

);

endmodule : cache
