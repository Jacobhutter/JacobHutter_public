library verilog;
use verilog.vl_types.all;
entity cache4 is
end cache4;
