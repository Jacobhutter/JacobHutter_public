library verilog;
use verilog.vl_types.all;
entity performence_counter_sv_unit is
end performence_counter_sv_unit;
