library verilog;
use verilog.vl_types.all;
entity MMIO_counter_sv_unit is
end MMIO_counter_sv_unit;
