library verilog;
use verilog.vl_types.all;
entity dirtywrite_sv_unit is
end dirtywrite_sv_unit;
