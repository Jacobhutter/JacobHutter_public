library verilog;
use verilog.vl_types.all;
entity cache4_datapath_sv_unit is
end cache4_datapath_sv_unit;
