library verilog;
use verilog.vl_types.all;
entity swapaddress4_sv_unit is
end swapaddress4_sv_unit;
