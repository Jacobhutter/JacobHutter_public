library verilog;
use verilog.vl_types.all;
entity datawrite_sv_unit is
end datawrite_sv_unit;
