import lc3b_types::*;

module cache_datapath
(
    input clk,


);

endmodule : cache_datapath
