library verilog;
use verilog.vl_types.all;
entity ebhitchecker_sv_unit is
end ebhitchecker_sv_unit;
