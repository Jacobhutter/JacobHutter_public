library verilog;
use verilog.vl_types.all;
entity exmem_sv_unit is
end exmem_sv_unit;
