library verilog;
use verilog.vl_types.all;
entity lruwrite_sv_unit is
end lruwrite_sv_unit;
