library verilog;
use verilog.vl_types.all;
entity dataforward_sv_unit is
end dataforward_sv_unit;
