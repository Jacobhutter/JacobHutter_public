library verilog;
use verilog.vl_types.all;
entity memwb_sv_unit is
end memwb_sv_unit;
