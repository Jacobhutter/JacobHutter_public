library verilog;
use verilog.vl_types.all;
entity selectway_sv_unit is
end selectway_sv_unit;
