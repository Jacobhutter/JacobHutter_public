library verilog;
use verilog.vl_types.all;
entity ebcontrol_sv_unit is
end ebcontrol_sv_unit;
