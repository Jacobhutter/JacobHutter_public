library verilog;
use verilog.vl_types.all;
entity ifid_sv_unit is
end ifid_sv_unit;
