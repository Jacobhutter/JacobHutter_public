library verilog;
use verilog.vl_types.all;
entity idex_sv_unit is
end idex_sv_unit;
