library verilog;
use verilog.vl_types.all;
entity global_bht_sv_unit is
end global_bht_sv_unit;
