module rowmodule( input Clk,Reset,

);


endmodule 
