import lc3b_types::*;

module cpu(
  instructions,
  data
);

cpu_datapath cd();

endmodule : cpu
